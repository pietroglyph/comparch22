`timescale 1ns / 100ps
`default_nettype none

`include "i2c_types.sv"

// TI has a good reference on how i2c works: https://training.ti.com/sites/default/files/docs/slides-i2c-protocol.pdf
// In this guide the "main" device is called the "controller" and the "secondary" device is called the "target".
module i2c_controller(
  clk, rst,
  scl, sda, mode,
  i_ready, i_valid, i_addr, i_data,
  o_ready, o_valid, o_data
);

parameter CLK_HZ = 12_000_000;
parameter I2C_CLK_HZ = 100_000; // Must be <= 400kHz
parameter DIVIDER_COUNT = CLK_HZ/I2C_CLK_HZ/2;  // Divide by two necessary since we toggle the signal
`ifdef SIMULATION
parameter COOLDOWN_CYCLES = 12; // Wait between transactions (can help smooth over issues with ACK or STOP or START conditions).
`else
parameter COOLDOWN_CYCLES = 120; // Wait between transactions (can help smooth over issues with ACK or STOP or START conditions).
`endif // SIMULATION

//Module I/O and parameters
input wire clk, rst; // standard signals
output logic scl; // i2c signals
inout wire sda;

// Create a tristate for the sda input/output pin.
// Tristates let you go into "high impedance" mode which allows the secondary device to use the same wire to send data back!
// It's your job to drive sda_oe (output enable) low (combinationally) when it's the secondary's turn to talk.
logic sda_oe; // output enable for the sda tristate
logic sda_out; // input to the tristate
assign sda = sda_oe ? sda_out : 1'bz; // Needs to be an assign, not always_comb for icarus verilog.

input wire i2c_transaction_t mode; // See i2c_types.sv, 0 is WRITE and 1 is READ
output logic i_ready; // ready/valid handshake signals
input wire i_valid;
input wire [6:0] i_addr; // the address of the secondary device.
input wire [7:0] i_data; // data to be sent on a WRITE opearation
input wire o_ready; // unused (for now)
output logic o_valid; // high when data is valid. Should stay high until a new i_valid starts a new transaction.
output logic [7:0] o_data; // the result of a read transaction (can be x's on a write).

// Main FSM logic
i2c_state_t state; // see i2c_types for the canonical states.

logic [$clog2(DIVIDER_COUNT):0] clk_divider_counter;
logic [$clog2(COOLDOWN_CYCLES):0] cooldown_counter; // optional, but recommended - have the system wait a few clk cycles before i_ready goes high again - this can make debugging STOP/ACK/START issues way easier!!!
logic [3:0] bit_counter;
logic [7:0] addr_buffer;
logic [7:0] data_buffer;

always_ff @(posedge clk) begin : i2c_fsm  
  if(rst) begin
    clk_divider_counter <= ($clog2(DIVIDER_COUNT)+1)'(DIVIDER_COUNT-1);
    cooldown_counter <= COOLDOWN_CYCLES;
    bit_counter <= 0;
    scl <= 1;
    o_data <= 0;
    o_valid <= 0;
    i_ready <= 1;
    state <= S_IDLE;
  end else begin // out of reset
	  if (state == S_IDLE) begin
		  // Reset SCL; it will be set low next state (i.e. after
		  // cooldown and one divided clock)
		  scl <= 1;
		  // Immediately enable setting SDA; we have a combinational
		  // logic block below that will then effectively pull SDA
		  // low.
		  if (i_valid & i_ready) begin
			  // We want the counter to be correct for when we
			  // return to S_IDLE.
			  cooldown_counter <= COOLDOWN_CYCLES;
			  // We want this counter to be correct when we
			  // transition to the next state.
			  clk_divider_counter <= ($clog2(DIVIDER_COUNT)+1)'(DIVIDER_COUNT-1);

			  // We need to sample the requested address and data
			  // to write (even if it may not be written) only
			  // when i_valid is true and when we're valid.
			  // Otherwise our "contract" with other modules is
			  // that we'll ignore those inputs.
			  addr_buffer <= {i_addr, mode};
			  data_buffer <= i_data;

			  // We're leaving idle, so the output is not going to
			  // be valid anymore.
			  o_valid <= 0;
			  // That also means that we're not ready to recieve
			  // input anymore, because we're going to be
			  // (potentially) writing whatever input data we were
			  // given.
			  i_ready <= 0;
			  state <= S_START;
		  end else if (~i_ready) begin
			  if (cooldown_counter == 0) i_ready <= 1;
			  else begin
				  i_ready <= 0;
				  cooldown_counter <= cooldown_counter - 1;
			  end
		  end
	  end else if (clk_divider_counter == 0) begin
		  clk_divider_counter <= ($clog2(DIVIDER_COUNT)+1)'(DIVIDER_COUNT-1);

		  scl <= ~scl;
		  case (state)
			  S_START: begin // All we do is bring scl low (see above), reset bit counter, and go next
				  state <= S_ADDR;
				  // We will write out 7 bits plus
				  // a read/write bit (i.e. addr_buffer's max
				  // index is 7). We start at the max index
				  // because we write the address out in
				  // little endian.
				  bit_counter <= 7;
			  end
			  S_ADDR: begin
				  // Only change the bit to write out on
				  // a negative edge.
				  if (scl) begin
					  if (bit_counter == 0) state <= S_ACK_ADDR;
					  else bit_counter <= bit_counter - 1;
				  end
			  end
			  S_ACK_ADDR: begin
				  `ifndef SIMULATION
				  if (~sda) begin
				  `endif
					  if (scl & addr_buffer[0] == WRITE_8BIT_REGISTER) state <= S_WR_DATA;
					  else if (~scl & addr_buffer[0] == READ_8BIT) state <= S_RD_DATA;
				  `ifndef SIMULATION
				  end
				  `endif

				  // We need to read or write 8 bits in the
				  // next state.
				  bit_counter <= 7;
			  end
			  S_WR_DATA: begin
				  // Only change the bit to write out on
				  // a negative edge.
				  if (scl) begin
					  if (bit_counter == 0) state <= S_ACK_WR;
					  else bit_counter <= bit_counter - 1;
				  end
			  end
			  S_ACK_WR: begin
				  // We want to transition on a rising edge,
				  // because we want SCL to be high first
				  // (before SDA goes high in stop).
				  if (~sda & scl) state <= S_STOP;
			  end
			  S_RD_DATA: begin
				  // Only change the bit to read on a positive
				  // edge (the secondary should be setting on
				  // a negative edge).
				  if (~scl) begin
					  data_buffer[bit_counter[2:0]] <= sda;
					  if (bit_counter == 0) state <= S_ACK_RD;
					  else bit_counter <= bit_counter - 1;
				  end
			  end
			  S_ACK_RD: begin
				  // SDA gets pulled low combinationally (see
				  // below).
				  
				  // We want to transition on a rising edge,
				  // because we want SCL to be high first
				  // (before SDA goes high in stop).
				  if (~scl) begin
					  state <= S_STOP;
					  // Target sent an ACK so the data we read
					  // should be good.
					  o_valid <= 1;
					  // Need to copy into data buffer.
					  o_data <= data_buffer;
				  end
			  end
			  S_STOP: begin
				  state <= S_IDLE;
			  end
			  default: state <= S_ERROR;
		  endcase
	  end else clk_divider_counter <= clk_divider_counter - 1;
  end
end

always_comb case (state)
	S_IDLE, S_START, S_ADDR, S_WR_DATA, S_ACK_RD, S_STOP: sda_oe = 1;
	default: sda_oe = 0;
endcase

always_comb case (state)
	S_IDLE: sda_out = 1;
	// We ensure SCL is high in start, so we pull SDA low to get the start
	// condition.
	S_START: sda_out = 0;
	S_ADDR: sda_out = addr_buffer[bit_counter[2:0]];
	// We go into this state immediately, but wait one divided clock cycle to
	// get to a case where we set sda_oe = 0.
	S_WR_DATA: sda_out = data_buffer[bit_counter[2:0]];
	S_ACK_RD: sda_out = 0;
	S_STOP: sda_out = 0;
	// We don't explicitly pull SDA up on idle (or stop??); instead, we set
	// the ouput to high impedence, and SDA gets pulled up. Other
	// controllers will detect the stop condition, and can trigger their
	// own start condition as soon as they want.
	default: sda_out = 0; // Doesn't matter, tri-state buffer is high impedance
endcase

endmodule
